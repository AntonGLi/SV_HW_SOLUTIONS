//
//  schoolRISCV - small RISC-V CPU
//
//  Originally based on Sarah L. Harris MIPS CPU
//  & schoolMIPS project.
//
//  Copyright (c) 2017-2020 Stanislav Zhelnio & Aleksandr Romanov.
//
//  Modified in 2024 by Yuri Panchul & Mike Kuskov
//  for systemverilog-homework project.
//

`include "sr_cpu.sv"

module srat_cpu
(
    input           clk,      // clock
    input           rst,      // reset

    output  [31:0]  imAddr,   // instruction memory address
    input   [31:0]  imData,   // instruction memory data

    input   [ 4:0]  regAddr,  // debug access reg address
    output  [31:0]  regData   // debug access reg data
);
    // control wires

    wire        aluZero;
    wire        pcSrc;
    wire        regWrite;
    wire        aluSrc;
    wire        wdSrc;
    wire  [2:0] aluControl;

    // instruction decode wires

    wire [ 6:0] cmdOp;
    wire [ 4:0] rd;
    wire [ 2:0] cmdF3;
    wire [ 4:0] rs1;
    wire [ 4:0] rs2;
    wire [ 6:0] cmdF7;
    wire [31:0] immI;
    wire [31:0] immB;
    wire [31:0] immU;
	 wire [31:0] IMM_J;
	 
	 wire [31:0] rd0;
    wire [31:0] rd1;
    wire [31:0] rd2;
    wire [31:0] wd3;
	 wire pc_JAL;

	 //MUL
	 wire [31:0] res_mul;
	   wire [31:0] pc;
	 
	 wire vld_mul;
	 wire start = (aluControl == `ALU_MUL);

	 wire [31:0] srcB = aluSrc ? immI :
								(pc_JAL) ? 32'd4 : rd2;
	 
	 wire [31:0] srcA = (pc_JAL) ? pc : rd1;
	 
    mul mul_11
    (
    .clk(clk),
    .rst(rst),

    .a(srcA),
    .b(srcB),

    .start(start) ,

    .res_mul(res_mul),
    .end_mul(vld_mul)
);

	 
    // program counter

    wire [31:0] pcBranch = pc + immB;
    wire [31:0] pcPlus4  = pc + 32'd4;
	 wire [31:0] pcJAL = pc + IMM_J;
    wire [31:0] pc_mul   = (vld_mul) ? (pc + 32'd4) : (pc);

    wire [31:0] pcNext   = (pc_JAL) ? pcJAL :
									(pcSrc) ? pcBranch :
									(aluControl == `ALU_MUL) ? pc_mul:
														           pcPlus4;

    register_with_rst r_pc (clk, rst, pcNext, pc);

    // program memory access

    assign imAddr = pc >> 2;
    wire [31:0] instr = imData;

    // instruction decode

    sr_decode id
    (
        .instr      ( instr       ),
        .cmdOp      ( cmdOp       ),
        .rd         ( rd          ),
        .cmdF3      ( cmdF3       ),
        .rs1        ( rs1         ),
        .rs2        ( rs2         ),
        .cmdF7      ( cmdF7       ),
        .immI       ( immI        ),
        .immB       ( immB        ),
        .immU       ( immU        ),
		  .IMM_J (IMM_J)
    );

    // register file



    sr_register_file i_rf
    (
        .clk        ( clk         ),
        .a0         ( regAddr     ),
        .a1         ( rs1         ),
        .a2         ( rs2         ),
        .a3         ( rd          ),
        .rd0        ( rd0         ),
        .rd1        ( rd1         ),
        .rd2        ( rd2         ),
        .wd3        ( wd3         ),
        .we3        ( regWrite    )
    );

    // alu


    wire [31:0] aluResult_nomul;
	 wire [31:0] aluResult;
	 assign aluResult = (vld_mul) ? res_mul : aluResult_nomul;

    sr_alu alu
    (
        .srcA       ( srcA         ),
        .srcB       ( srcB        ),
        .oper       ( aluControl  ),
        .zero       ( aluZero     ),
        .result     ( aluResult_nomul   )
    );

    assign wd3 = wdSrc ? immU : aluResult;

    // control

    sr_control sm_control
    (
        .cmdOp      ( cmdOp       ),
        .cmdF3      ( cmdF3       ),
        .cmdF7      ( cmdF7       ),
        .aluZero    ( aluZero     ),
        .pcSrc      ( pcSrc       ),
        .regWrite   ( regWrite    ),
        .aluSrc     ( aluSrc      ),
        .wdSrc      ( wdSrc       ),
        .aluControl ( aluControl  ),
		  .vld (vld_mul),
		  .pc_JAL (pc_JAL)

    );

    // debug register access

    assign regData = (regAddr != '0) ? rd0 : pc;

endmodule